module Execute(
    input wire clk, regdst, alusrc,
    input wire input_WB,
    input wire input_m,
    input wire instr_2016,
    output wire Latch_Mem
    );
    
endmodule